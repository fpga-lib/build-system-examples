//-------------------------------------------------------------------------------
//
//     Project: Any
//
//     Purpose: Adder module. Wraps HLS-generated module
//
//-------------------------------------------------------------------------------

`include "cfg_params.svh"

//-------------------------------------------------------------------------------
module automatic adder_m
(
    input logic  clk,
    input logic  rst,

    dinp_if.s    a,
    dinp_if.s    b,
    dout_if.m    out
);

//------------------------------------------------------------------------------
//
//    Settings
//
    
//------------------------------------------------------------------------------
//
//    Types
//


//------------------------------------------------------------------------------
//
//    Objects
//
logic ap_local_block;
logic ap_local_deadlock;

//------------------------------------------------------------------------------
//
//    Functions and tasks
//

//------------------------------------------------------------------------------
//
//    Logic
//

//------------------------------------------------------------------------------
//
//    Instances
//
adder_hlsip adder_hls
(
    .ap_clk            (  clk              ),
    .ap_rst            (  rst              ),
    .ap_local_block    ( ap_local_block    ),
    .ap_local_deadlock ( ap_local_deadlock ),
    .a_ap_vld          ( a.valid           ),
    .a                 ( a.data            ),
    .b_ap_vld          ( b.valid           ),
    .b                 ( b.data            ),
    .out_r_ap_vld      ( out.valid         ),
    .out_r             ( out.data          )
);
//-------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------

